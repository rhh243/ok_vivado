//------------------------------------------------------------------------
// okHostCallsSecondary.vh
//
// Description:
//    This file is included by a test fixture designed to mimic FrontPanel
//    operations.  The functions and task below provide a pseudo
//    translation between the FrontPanel operations and the hi_cmd, hi_out,
//    and hi_inout signals.
//
//    Note that this file is designed to mimic a secondary FrontPanel
//    interface. Use of this file assumes a primary FrontPanel interface
//    is used in the same simulation and that okHostCalls.v for the primary
//    interface is included prior to inclusion of this file.
//------------------------------------------------------------------------
// Copyright (c) 2022 Opal Kelly Incorporated
//------------------------------------------------------------------------

//------------------------------------------------------------------------
// *  Do not edit any of the defines, registers, integers, arrays, or
//    functions below this point.
// *  Tasks in Verilog cannot pass arrays.  The pipe tasks utilize arrays
//    of data. If you require multiple pipe arrays, you may create new
//    arrays in the top level file (that `includes this file), duplicate
//    the pipe tasks below as required, change the names of the duplicated
//    tasks to unique identifiers, and alter the pipe array in those tasks
//    to your newly generated arrays in the top level file.
// *  For example, in the top level file, along with:
//       reg   [7:0] pipeIn_s [0:(pipeInSize-1)];
//       reg   [7:0] pipeOut_s [0:(pipeOutSize-1)];
//       - Add:   reg   [7:0] pipeIn2_s [0:1023];
//       - Then, copy the WriteToPipeInSecondary task here, rename it
//         WriteToPipeInSecondary2, and finally change pipeIn_s[i] in
//         WriteToPipeInSecondary2 to pipeIn2_s[i].
//    The task and operation can then be called with a:
//       WriteToPipeInSecondary2(8'h80, 1024);//endpoint 0x80 pipe received pipeIn2_s
//------------------------------------------------------------------------
                 
// Local okHostCall signals
reg            hi_clk_s;
reg            hi_drive_s;
reg   [2:0]    hi_cmd_s;
wire           hi_busy_s;
wire  [31:0]   hi_datain_s;
reg   [31:0]   hi_dataout_s;

reg   [31:0]   WireIns_s [0:31];   // 32x32 array storing WireIn values
reg   [31:0]   WireOuts_s [0:31];  // 32x32 array storing WireOut values
reg   [31:0]   Triggered_s [0:31]; // 32x32 array storing IsTriggered values

initial begin
	hi_clk_s     = 1'b0;
	hi_drive_s   = 1'b0;
	hi_cmd_s     = `DNOP;
	hi_dataout_s = 32'h0000;
end

// Mapping of local okHostCall signals to okHost interface
assign okUHs[0]   = hi_clk_s;
assign okUHs[1]   = hi_drive_s;
assign okUHs[4:2] = hi_cmd_s; 
assign hi_datain_s = okUHUs;
assign hi_busy_s   = okHUs[0]; 
assign okUHUs     = hi_drive_s ? hi_dataout_s : 32'hzzzz;

// Clock Generation
always #tCK hi_clk_s = ~hi_clk_s;
	
//---------------------------------------------------------
// FrontPanelReset
//---------------------------------------------------------
task FrontPanelResetSecondary ();
	integer i;
begin
	for (i=0; i<32; i=i+1) begin
		WireIns_s[i] = 32'h0000;
		WireOuts_s[i] = 32'h0000;
		Triggered_s[i] = 32'h0000;
	end
	
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DReset;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DNOP;
	wait (hi_busy_s == 0);
end
endtask

//---------------------------------------------------------
// SetWireInValue
//---------------------------------------------------------
task SetWireInValueSecondary (
	input    [7:0]    ep,
	input    [31:0]   val,
	input    [31:0]   mask
);
	reg   [31:0]   tmp;
begin
	tmp = WireIns_s[ep] & ~mask;
	WireIns_s[ep] = tmp | (val & mask);
end
endtask

//---------------------------------------------------------
// GetWireOutValue
//---------------------------------------------------------
function [31:0] GetWireOutValueSecondary (
	input    [7:0]    ep
);
begin
	GetWireOutValueSecondary = WireOuts_s[ep - 8'h20];
end
endfunction

//---------------------------------------------------------
// IsTriggered
//---------------------------------------------------------
function IsTriggeredSecondary (
	input    [7:0]    ep,
	input    [31:0]   mask
);
begin
	if ((Triggered_s[ep - 8'h60] & mask) >= 0) begin
		if ((Triggered_s[ep - 8'h60] & mask) == 0) begin
			IsTriggeredSecondary = 0;
		end else begin
			IsTriggeredSecondary = 1;
		end
	end else begin
		$display("***FRONTPANEL ERROR: IsTriggered Secondary mask 0x%04h covers unused Triggers", mask);
		IsTriggeredSecondary = 0;
	end
end
endfunction

//---------------------------------------------------------
// UpdateWireIns
//---------------------------------------------------------
task UpdateWireInsSecondary ();
   integer i;
begin
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DWires;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DUpdateWireIns;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DNOP;
	for (i=0; i<32; i=i+1) begin
		hi_dataout_s = WireIns_s[i];
		@(posedge hi_clk_s) ;
	end
	wait (hi_busy_s == 0);
end
endtask

//---------------------------------------------------------
// UpdateWireOuts
//---------------------------------------------------------
task UpdateWireOutsSecondary ();
	integer i;
begin
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DWires;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DUpdateWireOuts;
	@(posedge hi_clk_s);
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DNOP;
	@(posedge hi_clk_s) hi_drive_s = 0;
	@(posedge hi_clk_s); @(posedge hi_clk_s);
	for (i=0; i<32; i=i+1)
		@(posedge hi_clk_s) WireOuts_s[i] = hi_datain_s;
	wait (hi_busy_s == 0);
end
endtask

//---------------------------------------------------------
// ActivateTriggerIn
//---------------------------------------------------------
task ActivateTriggerInSecondary (
	input    [7:0]    ep,
	input    [31:0]  trig_bit
);
begin
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DTriggers;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DActivateTriggerIn;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_dataout_s = {24'h00, ep};
	@(posedge hi_clk_s) hi_dataout_s = (1'b1 << trig_bit);
	hi_cmd_s[2:0] = `DNOP;
	@(posedge hi_clk_s) hi_dataout_s = 32'h0000;
	wait (hi_busy_s == 0);
end
endtask

//---------------------------------------------------------
// UpdateTriggerOuts
//---------------------------------------------------------
task UpdateTriggerOutsSecondary ();
	integer i;
begin
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DTriggers;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DUpdateTriggerOuts;
	@(posedge hi_clk_s);
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DNOP;
	@(posedge hi_clk_s) hi_drive_s = 0;
	@(posedge hi_clk_s); @(posedge hi_clk_s); @(posedge hi_clk_s);
	
	for (i=0; i<UPDATE_TO_READOUT_CLOCKS; i=i+1)@(posedge hi_clk_s);
	
	for (i=0; i<32; i=i+1)
		@(posedge hi_clk_s) Triggered_s[i] = hi_datain_s;
	wait (hi_busy_s == 0);
end
endtask


//---------------------------------------------------------
// WriteToPipeIn
//---------------------------------------------------------
task WriteToPipeInSecondary (
	input    [7:0]    ep,
	input    [31:0]   length
);
	integer  len, i, j, k, blockSize;
begin
	len = length/4; j = 0; blockSize = 1024;
	if (length%2)
		$display("Error. Pipes commands may only send and receive an even # of bytes.");
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DPipes;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DWriteToPipeIn;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_dataout_s = {BlockDelayStates, ep};
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DNOP;
	hi_dataout_s = len;
	for (i=0; i < length; i=i+4) begin
		@(posedge hi_clk_s);
		hi_dataout_s[7:0]   = pipeIn_s[i];
		hi_dataout_s[15:8]  = pipeIn_s[i+1];
		hi_dataout_s[23:16] = pipeIn_s[i+2];
		hi_dataout_s[31:24] = pipeIn_s[i+3];
		j=j+4;
		if (j == blockSize) begin
			for (k=0; k < BlockDelayStates; k=k+1) begin
				@(posedge hi_clk_s);
			end
			j=0;
		end
	end
	wait (hi_busy_s == 0);
end
endtask


//---------------------------------------------------------
// ReadFromPipeOut
//---------------------------------------------------------
task ReadFromPipeOutSecondary (
	input    [7:0]    ep,
	input    [31:0]   length
);
	integer len, i, j, k, blockSize;
begin
	len = length/4; j = 0; blockSize = 1024;
	if (length%2)
		$display("Error. Pipes commands may only send and receive an even # of bytes.");
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DPipes;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DReadFromPipeOut;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_dataout_s = {BlockDelayStates, ep};
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DNOP;
	hi_dataout_s = len;
	@(posedge hi_clk_s) hi_drive_s = 0;
	for (i=0; i < length; i=i+4) begin
		@(posedge hi_clk_s);
		pipeOut_s[i]   = hi_datain_s[7:0];
		pipeOut_s[i+1] = hi_datain_s[15:8];
		pipeOut_s[i+2] = hi_datain_s[23:16];
		pipeOut_s[i+3] = hi_datain_s[31:24];
		j=j+4;
		if (j == blockSize) begin
			for (k=0; k < BlockDelayStates; k=k+1) begin
				@(posedge hi_clk_s);
			end
			j=0;
		end
	end
	wait (hi_busy_s == 0);
end
endtask

//---------------------------------------------------------
// WriteToBlockPipeIn
//---------------------------------------------------------
task WriteToBlockPipeInSecondary (
	input    [7:0]    ep,
	input    [31:0]   blockLength,
	input    [31:0]   length
);
	integer len, blockSize, blockNum, i, j, k;
begin
	len = length/4; blockSize = blockLength/4; k = 0;
	blockNum = len/blockSize;
	if (length%2)
		$display("Error. Pipes commands may only send and receive an even # of bytes.");
	if (blockLength%2)
		$display("Error. Block Length may only be an even # of bytes.");
	if (length%blockLength)
		$display("Error. Pipe length MUST be a multiple of block length!");
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DPipes;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DWriteToBlockPipeIn;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_dataout_s = {BlockDelayStates, ep};
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DNOP;
	hi_dataout_s = len;
	@(posedge hi_clk_s) hi_dataout_s = blockSize;
	@(posedge hi_clk_s) hi_dataout_s[7:0] = ReadyCheckDelay; hi_dataout_s[15:8] = PostReadyDelay;
	for (i=0; i < blockNum; i=i+1) begin
		while (hi_busy_s === 1) @(posedge hi_clk_s);
		while (hi_busy_s === 0) @(posedge hi_clk_s);
		@(posedge hi_clk_s); @(posedge hi_clk_s);
		for (j=0; j<blockSize; j=j+1) begin
			hi_dataout_s[7:0]   = pipeIn_s[k]; 
			hi_dataout_s[15:8]  = pipeIn_s[k+1];
			hi_dataout_s[23:16] = pipeIn_s[k+2];
			hi_dataout_s[31:24] = pipeIn_s[k+3];
			@(posedge hi_clk_s); k=k+4;
		end
		for (j=0; j < BlockDelayStates; j=j+1) @(posedge hi_clk_s);
	end
	wait (hi_busy_s == 0);
end
endtask

//---------------------------------------------------------
// ReadFromBlockPipeOut
//---------------------------------------------------------
task ReadFromBlockPipeOutSecondary (
	input    [7:0]    ep,
	input    [31:0]   blockLength,
	input    [31:0]   length
);
   integer len, blockSize, blockNum, i, j, k;
begin
	len = length/4; blockSize = blockLength/4; k = 0;
	blockNum = len/blockSize;
	if (length%2)
		$display("Error. Pipes commands may only send and receive an even # of bytes.");
	if (blockLength%2)
		$display("Error. Block Length may only be an even # of bytes.");
	if (length%blockLength)
		$display("Error. Pipe length MUST be a multiple of block length!");
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DPipes;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DReadFromBlockPipeOut;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_dataout_s = {BlockDelayStates, ep};
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DNOP;
	hi_dataout_s = len;
	@(posedge hi_clk_s) hi_dataout_s = blockSize;
	@(posedge hi_clk_s) hi_dataout_s[7:0] = ReadyCheckDelay; hi_dataout_s[15:8] = PostReadyDelay;
	@(posedge hi_clk_s) hi_drive_s = 0;
	for (i=0; i < blockNum; i=i+1) begin
		while (hi_busy_s === 1) @(posedge hi_clk_s);
		while (hi_busy_s === 0) @(posedge hi_clk_s);
		@(posedge hi_clk_s); @(posedge hi_clk_s);
		for (j=0; j<blockSize; j=j+1) begin
			pipeOut_s[k]   = hi_datain_s[7:0]; 
			pipeOut_s[k+1] = hi_datain_s[15:8];
			pipeOut_s[k+2] = hi_datain_s[23:16];
			pipeOut_s[k+3] = hi_datain_s[31:24];
			@(posedge hi_clk_s) k=k+4;
		end
		for (j=0; j < BlockDelayStates; j=j+1) @(posedge hi_clk_s);
	end
	wait (hi_busy_s == 0);
end
endtask

//---------------------------------------------------------
// WriteRegister
//---------------------------------------------------------
task WriteRegisterSecondary (
	input    [31:0]   address,
	input    [31:0]   data
);
begin
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DRegisters;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DWriteRegister;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_cmd_s[2:0] = `DNOP;
	@(posedge hi_clk_s) hi_dataout_s = address;
	@(posedge hi_clk_s) hi_dataout_s = data;
	wait (hi_busy_s == 0); hi_drive_s = 0; 
end
endtask

//---------------------------------------------------------
// ReadRegister
//---------------------------------------------------------
task ReadRegisterSecondary (
	input    [31:0]   address,
	output   [31:0]   data
);
begin
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DRegisters;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DReadRegister;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_cmd_s[2:0] = `DNOP;
	@(posedge hi_clk_s) hi_dataout_s = address;
	@(posedge hi_clk_s); hi_drive_s = 0; 
	@(posedge hi_clk_s);
	@(posedge hi_clk_s) data = hi_datain_s;
	wait (hi_busy_s == 0);
end
endtask

//---------------------------------------------------------
// WriteRegisterSet
//---------------------------------------------------------
task WriteRegisterSetSecondary ();
	integer i;
begin
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DRegisters;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DWriteRegisterSet;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_cmd_s[2:0] = `DNOP;
	@(posedge hi_clk_s); hi_dataout_s = u32Count_s;
	for (i=0; i < u32Count_s; i=i+1) begin
		@(posedge hi_clk_s) hi_dataout_s = u32Address_s[i];
		@(posedge hi_clk_s) hi_dataout_s = u32Data_s[i];
		@(posedge hi_clk_s); @(posedge hi_clk_s); 
	end
	wait (hi_busy_s == 0); hi_drive_s = 0; 
end
endtask

//---------------------------------------------------------
// ReadRegisterSet
//---------------------------------------------------------
task ReadRegisterSetSecondary ();
	integer i;
begin
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DRegisters;
	@(posedge hi_clk_s) hi_cmd_s[2:0] = `DReadRegisterSet;
	@(posedge hi_clk_s);
	hi_drive_s = 1;
	hi_cmd_s[2:0] = `DNOP;
	@(posedge hi_clk_s); hi_dataout_s = u32Count_s;
	for (i=0; i < u32Count_s; i=i+1) begin
		@(posedge hi_clk_s) hi_dataout_s = u32Address_s[i];
		@(posedge hi_clk_s); hi_drive_s = 0; 
		@(posedge hi_clk_s);
		@(posedge hi_clk_s) u32Data_s[i] = hi_datain_s;
		hi_drive_s = 1;
	end
	wait (hi_busy_s == 0);
end
endtask
